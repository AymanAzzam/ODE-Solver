/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed Apr 22 04:57:20 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2696149395 */

module Add_Sub(A, B, result, overflow);
   input [15:0]A;
   input [15:0]B;
   output [15:0]result;
   output overflow;

   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;

   XOR2_X1 i_0_0_0 (.A(A[0]), .B(B[0]), .Z(result[0]));
   XNOR2_X1 i_0_0_1 (.A(n_0_0_5), .B(n_0_0_0), .ZN(result[1]));
   NOR2_X1 i_0_0_2 (.A1(n_0_0_58), .A2(n_0_0_6), .ZN(n_0_0_0));
   XNOR2_X1 i_0_0_3 (.A(n_0_0_4), .B(n_0_0_1), .ZN(result[2]));
   XNOR2_X1 i_0_0_4 (.A(A[2]), .B(B[2]), .ZN(n_0_0_1));
   XNOR2_X1 i_0_0_5 (.A(n_0_0_7), .B(n_0_0_2), .ZN(result[3]));
   NAND2_X1 i_0_0_6 (.A1(n_0_0_60), .A2(n_0_0_3), .ZN(n_0_0_2));
   OAI21_X1 i_0_0_7 (.A(n_0_0_4), .B1(B[2]), .B2(A[2]), .ZN(n_0_0_3));
   OAI21_X1 i_0_0_8 (.A(n_0_0_59), .B1(n_0_0_6), .B2(n_0_0_5), .ZN(n_0_0_4));
   NAND2_X1 i_0_0_9 (.A1(A[0]), .A2(B[0]), .ZN(n_0_0_5));
   NOR2_X1 i_0_0_10 (.A1(A[1]), .A2(B[1]), .ZN(n_0_0_6));
   XNOR2_X1 i_0_0_11 (.A(A[3]), .B(B[3]), .ZN(n_0_0_7));
   XOR2_X1 i_0_0_12 (.A(n_0_0_55), .B(n_0_0_51), .Z(result[4]));
   XNOR2_X1 i_0_0_13 (.A(n_0_0_13), .B(n_0_0_8), .ZN(result[5]));
   XNOR2_X1 i_0_0_14 (.A(A[5]), .B(B[5]), .ZN(n_0_0_8));
   XNOR2_X1 i_0_0_15 (.A(n_0_0_11), .B(n_0_0_9), .ZN(result[6]));
   XOR2_X1 i_0_0_16 (.A(A[6]), .B(B[6]), .Z(n_0_0_9));
   XNOR2_X1 i_0_0_17 (.A(n_0_0_14), .B(n_0_0_10), .ZN(result[7]));
   OAI21_X1 i_0_0_18 (.A(n_0_0_49), .B1(n_0_0_11), .B2(n_0_0_62), .ZN(n_0_0_10));
   OR2_X1 i_0_0_19 (.A1(n_0_0_54), .A2(n_0_0_12), .ZN(n_0_0_11));
   AOI21_X1 i_0_0_20 (.A(n_0_0_13), .B1(B[5]), .B2(A[5]), .ZN(n_0_0_12));
   OAI21_X1 i_0_0_21 (.A(n_0_0_52), .B1(n_0_0_53), .B2(n_0_0_55), .ZN(n_0_0_13));
   NAND2_X1 i_0_0_22 (.A1(n_0_0_47), .A2(n_0_0_45), .ZN(n_0_0_14));
   NOR2_X1 i_0_0_23 (.A1(n_0_0_43), .A2(n_0_0_15), .ZN(result[8]));
   AOI21_X1 i_0_0_24 (.A(n_0_0_44), .B1(n_0_0_45), .B2(n_0_0_46), .ZN(n_0_0_15));
   XNOR2_X1 i_0_0_25 (.A(n_0_0_21), .B(n_0_0_16), .ZN(result[9]));
   XOR2_X1 i_0_0_26 (.A(A[9]), .B(B[9]), .Z(n_0_0_16));
   XNOR2_X1 i_0_0_27 (.A(n_0_0_20), .B(n_0_0_17), .ZN(result[10]));
   XNOR2_X1 i_0_0_28 (.A(A[10]), .B(B[10]), .ZN(n_0_0_17));
   XNOR2_X1 i_0_0_29 (.A(n_0_0_22), .B(n_0_0_18), .ZN(result[11]));
   AOI21_X1 i_0_0_30 (.A(n_0_0_19), .B1(B[10]), .B2(A[10]), .ZN(n_0_0_18));
   AOI21_X1 i_0_0_31 (.A(n_0_0_40), .B1(n_0_0_21), .B2(n_0_0_63), .ZN(n_0_0_19));
   OAI21_X1 i_0_0_32 (.A(n_0_0_63), .B1(n_0_0_41), .B2(n_0_0_21), .ZN(n_0_0_20));
   AOI21_X1 i_0_0_33 (.A(n_0_0_43), .B1(B[8]), .B2(A[8]), .ZN(n_0_0_21));
   XOR2_X1 i_0_0_34 (.A(A[11]), .B(B[11]), .Z(n_0_0_22));
   XNOR2_X1 i_0_0_35 (.A(n_0_0_37), .B(n_0_0_23), .ZN(result[12]));
   XNOR2_X1 i_0_0_36 (.A(A[12]), .B(B[12]), .ZN(n_0_0_23));
   AND2_X1 i_0_0_37 (.A1(n_0_0_25), .A2(n_0_0_24), .ZN(result[13]));
   OAI21_X1 i_0_0_38 (.A(n_0_0_33), .B1(n_0_0_34), .B2(n_0_0_65), .ZN(n_0_0_24));
   NAND2_X1 i_0_0_39 (.A1(n_0_0_66), .A2(n_0_0_34), .ZN(n_0_0_25));
   XNOR2_X1 i_0_0_40 (.A(n_0_0_33), .B(n_0_0_26), .ZN(result[14]));
   XNOR2_X1 i_0_0_41 (.A(A[14]), .B(B[14]), .ZN(n_0_0_26));
   XNOR2_X1 i_0_0_42 (.A(n_0_0_30), .B(n_0_0_27), .ZN(result[15]));
   NOR2_X1 i_0_0_43 (.A1(n_0_0_29), .A2(n_0_0_28), .ZN(n_0_0_27));
   MUX2_X1 i_0_0_44 (.A(n_0_0_28), .B(n_0_0_29), .S(n_0_0_30), .Z(overflow));
   NOR2_X1 i_0_0_45 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0_28));
   AND2_X1 i_0_0_46 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0_29));
   AOI21_X1 i_0_0_47 (.A(n_0_0_31), .B1(B[14]), .B2(A[14]), .ZN(n_0_0_30));
   INV_X1 i_0_0_48 (.A(n_0_0_32), .ZN(n_0_0_31));
   OAI21_X1 i_0_0_49 (.A(n_0_0_33), .B1(B[14]), .B2(A[14]), .ZN(n_0_0_32));
   OAI21_X1 i_0_0_50 (.A(n_0_0_65), .B1(n_0_0_34), .B2(n_0_0_66), .ZN(n_0_0_33));
   AOI21_X1 i_0_0_51 (.A(n_0_0_35), .B1(B[12]), .B2(A[12]), .ZN(n_0_0_34));
   INV_X1 i_0_0_52 (.A(n_0_0_36), .ZN(n_0_0_35));
   OAI21_X1 i_0_0_53 (.A(n_0_0_37), .B1(B[12]), .B2(A[12]), .ZN(n_0_0_36));
   NOR2_X1 i_0_0_54 (.A1(n_0_0_64), .A2(n_0_0_38), .ZN(n_0_0_37));
   AOI221_X1 i_0_0_55 (.A(n_0_0_39), .B1(B[10]), .B2(A[10]), .C1(A[11]), 
      .C2(B[11]), .ZN(n_0_0_38));
   NOR2_X1 i_0_0_56 (.A1(n_0_0_42), .A2(n_0_0_40), .ZN(n_0_0_39));
   OAI22_X1 i_0_0_57 (.A1(A[10]), .A2(B[10]), .B1(B[9]), .B2(A[9]), .ZN(n_0_0_40));
   NOR2_X1 i_0_0_58 (.A1(A[9]), .A2(B[9]), .ZN(n_0_0_41));
   AOI21_X1 i_0_0_59 (.A(n_0_0_43), .B1(B[9]), .B2(A[9]), .ZN(n_0_0_42));
   AND3_X1 i_0_0_60 (.A1(n_0_0_46), .A2(n_0_0_45), .A3(n_0_0_44), .ZN(n_0_0_43));
   XOR2_X1 i_0_0_61 (.A(A[8]), .B(B[8]), .Z(n_0_0_44));
   OR2_X1 i_0_0_62 (.A1(A[7]), .A2(B[7]), .ZN(n_0_0_45));
   OAI21_X1 i_0_0_63 (.A(n_0_0_47), .B1(n_0_0_48), .B2(n_0_0_62), .ZN(n_0_0_46));
   NAND2_X1 i_0_0_64 (.A1(A[7]), .A2(B[7]), .ZN(n_0_0_47));
   AOI221_X1 i_0_0_65 (.A(n_0_0_50), .B1(B[5]), .B2(A[5]), .C1(A[6]), .C2(B[6]), 
      .ZN(n_0_0_48));
   NAND2_X1 i_0_0_66 (.A1(A[6]), .A2(B[6]), .ZN(n_0_0_49));
   NOR3_X1 i_0_0_67 (.A1(n_0_0_55), .A2(n_0_0_54), .A3(n_0_0_51), .ZN(n_0_0_50));
   XNOR2_X1 i_0_0_68 (.A(A[4]), .B(B[4]), .ZN(n_0_0_51));
   NAND2_X1 i_0_0_69 (.A1(A[4]), .A2(B[4]), .ZN(n_0_0_52));
   NOR2_X1 i_0_0_70 (.A1(A[4]), .A2(B[4]), .ZN(n_0_0_53));
   NOR2_X1 i_0_0_71 (.A1(A[5]), .A2(B[5]), .ZN(n_0_0_54));
   OAI21_X1 i_0_0_72 (.A(n_0_0_56), .B1(B[3]), .B2(A[3]), .ZN(n_0_0_55));
   NAND3_X1 i_0_0_73 (.A1(n_0_0_61), .A2(n_0_0_60), .A3(n_0_0_57), .ZN(n_0_0_56));
   OAI21_X1 i_0_0_74 (.A(n_0_0_58), .B1(B[2]), .B2(A[2]), .ZN(n_0_0_57));
   INV_X1 i_0_0_75 (.A(n_0_0_59), .ZN(n_0_0_58));
   NAND2_X1 i_0_0_76 (.A1(A[1]), .A2(B[1]), .ZN(n_0_0_59));
   NAND2_X1 i_0_0_77 (.A1(A[2]), .A2(B[2]), .ZN(n_0_0_60));
   NAND2_X1 i_0_0_78 (.A1(A[3]), .A2(B[3]), .ZN(n_0_0_61));
   NOR2_X1 i_0_0_79 (.A1(A[6]), .A2(B[6]), .ZN(n_0_0_62));
   NAND2_X1 i_0_0_80 (.A1(A[9]), .A2(B[9]), .ZN(n_0_0_63));
   NOR2_X1 i_0_0_81 (.A1(A[11]), .A2(B[11]), .ZN(n_0_0_64));
   NAND2_X1 i_0_0_82 (.A1(A[13]), .A2(B[13]), .ZN(n_0_0_65));
   NOR2_X1 i_0_0_83 (.A1(A[13]), .A2(B[13]), .ZN(n_0_0_66));
endmodule
