/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed Apr 22 04:59:39 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 618056553 */

module Add_Sub(A, B, result, overflow);
   input [15:0]A;
   input [15:0]B;
   output [15:0]result;
   output overflow;

   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;

   OAI33_X1 i_0_0_0 (.A1(n_0_0_55), .A2(n_0_0_9), .A3(n_0_0_62), .B1(A[15]), 
      .B2(n_0_0_8), .B3(B[15]), .ZN(overflow));
   AOI21_X1 i_0_0_1 (.A(n_0_0_31), .B1(n_0_0_56), .B2(n_0_0_49), .ZN(result[0]));
   XNOR2_X1 i_0_0_2 (.A(n_0_0_31), .B(n_0_0_0), .ZN(result[1]));
   OAI22_X1 i_0_0_3 (.A1(n_0_0_57), .A2(n_0_0_50), .B1(B[1]), .B2(A[1]), 
      .ZN(n_0_0_0));
   XNOR2_X1 i_0_0_4 (.A(n_0_0_32), .B(n_0_0_29), .ZN(result[2]));
   XNOR2_X1 i_0_0_5 (.A(n_0_0_27), .B(n_0_0_1), .ZN(result[3]));
   AOI22_X1 i_0_0_6 (.A1(n_0_0_58), .A2(A[3]), .B1(B[3]), .B2(n_0_0_51), 
      .ZN(n_0_0_1));
   XOR2_X1 i_0_0_7 (.A(n_0_0_25), .B(n_0_0_2), .Z(result[4]));
   AOI22_X1 i_0_0_8 (.A1(n_0_0_59), .A2(n_0_0_52), .B1(B[4]), .B2(A[4]), 
      .ZN(n_0_0_2));
   XNOR2_X1 i_0_0_9 (.A(n_0_0_23), .B(n_0_0_3), .ZN(result[5]));
   OAI22_X1 i_0_0_10 (.A1(n_0_0_60), .A2(n_0_0_53), .B1(B[5]), .B2(A[5]), 
      .ZN(n_0_0_3));
   XNOR2_X1 i_0_0_11 (.A(n_0_0_35), .B(n_0_0_21), .ZN(result[6]));
   XOR2_X1 i_0_0_12 (.A(n_0_0_20), .B(n_0_0_4), .Z(result[7]));
   OAI21_X1 i_0_0_13 (.A(n_0_0_37), .B1(B[7]), .B2(A[7]), .ZN(n_0_0_4));
   XNOR2_X1 i_0_0_14 (.A(n_0_0_39), .B(n_0_0_19), .ZN(result[8]));
   XOR2_X1 i_0_0_15 (.A(n_0_0_18), .B(n_0_0_5), .Z(result[9]));
   OAI21_X1 i_0_0_16 (.A(n_0_0_40), .B1(B[9]), .B2(A[9]), .ZN(n_0_0_5));
   XOR2_X1 i_0_0_17 (.A(n_0_0_41), .B(n_0_0_16), .Z(result[10]));
   XNOR2_X1 i_0_0_18 (.A(n_0_0_15), .B(n_0_0_6), .ZN(result[11]));
   OAI22_X1 i_0_0_19 (.A1(n_0_0_61), .A2(n_0_0_54), .B1(B[11]), .B2(A[11]), 
      .ZN(n_0_0_6));
   XNOR2_X1 i_0_0_20 (.A(n_0_0_44), .B(n_0_0_13), .ZN(result[12]));
   XOR2_X1 i_0_0_21 (.A(n_0_0_12), .B(n_0_0_7), .Z(result[13]));
   OAI21_X1 i_0_0_22 (.A(n_0_0_45), .B1(B[13]), .B2(A[13]), .ZN(n_0_0_7));
   XOR2_X1 i_0_0_23 (.A(n_0_0_46), .B(n_0_0_10), .Z(result[14]));
   XNOR2_X1 i_0_0_24 (.A(n_0_0_48), .B(n_0_0_9), .ZN(result[15]));
   INV_X1 i_0_0_25 (.A(n_0_0_9), .ZN(n_0_0_8));
   OAI21_X1 i_0_0_26 (.A(n_0_0_47), .B1(n_0_0_46), .B2(n_0_0_10), .ZN(n_0_0_9));
   OAI21_X1 i_0_0_27 (.A(n_0_0_11), .B1(B[13]), .B2(A[13]), .ZN(n_0_0_10));
   NAND2_X1 i_0_0_28 (.A1(n_0_0_45), .A2(n_0_0_12), .ZN(n_0_0_11));
   AOI22_X1 i_0_0_29 (.A1(B[12]), .A2(A[12]), .B1(n_0_0_43), .B2(n_0_0_13), 
      .ZN(n_0_0_12));
   AOI21_X1 i_0_0_30 (.A(n_0_0_14), .B1(n_0_0_61), .B2(n_0_0_54), .ZN(n_0_0_13));
   AOI21_X1 i_0_0_31 (.A(n_0_0_15), .B1(B[11]), .B2(A[11]), .ZN(n_0_0_14));
   OAI21_X1 i_0_0_32 (.A(n_0_0_42), .B1(n_0_0_41), .B2(n_0_0_16), .ZN(n_0_0_15));
   OAI21_X1 i_0_0_33 (.A(n_0_0_17), .B1(B[9]), .B2(A[9]), .ZN(n_0_0_16));
   NAND2_X1 i_0_0_34 (.A1(n_0_0_40), .A2(n_0_0_18), .ZN(n_0_0_17));
   AOI22_X1 i_0_0_35 (.A1(B[8]), .A2(A[8]), .B1(n_0_0_38), .B2(n_0_0_19), 
      .ZN(n_0_0_18));
   AOI21_X1 i_0_0_36 (.A(n_0_0_36), .B1(n_0_0_37), .B2(n_0_0_20), .ZN(n_0_0_19));
   AOI22_X1 i_0_0_37 (.A1(B[6]), .A2(A[6]), .B1(n_0_0_34), .B2(n_0_0_21), 
      .ZN(n_0_0_20));
   AOI21_X1 i_0_0_38 (.A(n_0_0_22), .B1(n_0_0_60), .B2(n_0_0_53), .ZN(n_0_0_21));
   AOI21_X1 i_0_0_39 (.A(n_0_0_23), .B1(B[5]), .B2(A[5]), .ZN(n_0_0_22));
   OAI21_X1 i_0_0_40 (.A(n_0_0_24), .B1(n_0_0_59), .B2(n_0_0_52), .ZN(n_0_0_23));
   OAI21_X1 i_0_0_41 (.A(n_0_0_25), .B1(B[4]), .B2(A[4]), .ZN(n_0_0_24));
   AOI21_X1 i_0_0_42 (.A(n_0_0_26), .B1(n_0_0_58), .B2(n_0_0_51), .ZN(n_0_0_25));
   AOI21_X1 i_0_0_43 (.A(n_0_0_27), .B1(B[3]), .B2(A[3]), .ZN(n_0_0_26));
   OAI21_X1 i_0_0_44 (.A(n_0_0_33), .B1(n_0_0_32), .B2(n_0_0_28), .ZN(n_0_0_27));
   INV_X1 i_0_0_45 (.A(n_0_0_29), .ZN(n_0_0_28));
   AOI21_X1 i_0_0_46 (.A(n_0_0_30), .B1(n_0_0_57), .B2(n_0_0_50), .ZN(n_0_0_29));
   AOI21_X1 i_0_0_47 (.A(n_0_0_31), .B1(B[1]), .B2(A[1]), .ZN(n_0_0_30));
   NOR2_X1 i_0_0_48 (.A1(n_0_0_56), .A2(n_0_0_49), .ZN(n_0_0_31));
   OAI21_X1 i_0_0_49 (.A(n_0_0_33), .B1(B[2]), .B2(A[2]), .ZN(n_0_0_32));
   NAND2_X1 i_0_0_50 (.A1(B[2]), .A2(A[2]), .ZN(n_0_0_33));
   INV_X1 i_0_0_51 (.A(n_0_0_35), .ZN(n_0_0_34));
   XNOR2_X1 i_0_0_52 (.A(B[6]), .B(A[6]), .ZN(n_0_0_35));
   NOR2_X1 i_0_0_53 (.A1(B[7]), .A2(A[7]), .ZN(n_0_0_36));
   NAND2_X1 i_0_0_54 (.A1(B[7]), .A2(A[7]), .ZN(n_0_0_37));
   INV_X1 i_0_0_55 (.A(n_0_0_39), .ZN(n_0_0_38));
   XNOR2_X1 i_0_0_56 (.A(B[8]), .B(A[8]), .ZN(n_0_0_39));
   NAND2_X1 i_0_0_57 (.A1(B[9]), .A2(A[9]), .ZN(n_0_0_40));
   OAI21_X1 i_0_0_58 (.A(n_0_0_42), .B1(B[10]), .B2(A[10]), .ZN(n_0_0_41));
   NAND2_X1 i_0_0_59 (.A1(B[10]), .A2(A[10]), .ZN(n_0_0_42));
   INV_X1 i_0_0_60 (.A(n_0_0_44), .ZN(n_0_0_43));
   XNOR2_X1 i_0_0_61 (.A(B[12]), .B(A[12]), .ZN(n_0_0_44));
   NAND2_X1 i_0_0_62 (.A1(B[13]), .A2(A[13]), .ZN(n_0_0_45));
   OAI21_X1 i_0_0_63 (.A(n_0_0_47), .B1(B[14]), .B2(A[14]), .ZN(n_0_0_46));
   NAND2_X1 i_0_0_64 (.A1(B[14]), .A2(A[14]), .ZN(n_0_0_47));
   AOI22_X1 i_0_0_65 (.A1(n_0_0_62), .A2(A[15]), .B1(B[15]), .B2(n_0_0_55), 
      .ZN(n_0_0_48));
   INV_X1 i_0_0_66 (.A(A[0]), .ZN(n_0_0_49));
   INV_X1 i_0_0_67 (.A(A[1]), .ZN(n_0_0_50));
   INV_X1 i_0_0_68 (.A(A[3]), .ZN(n_0_0_51));
   INV_X1 i_0_0_69 (.A(A[4]), .ZN(n_0_0_52));
   INV_X1 i_0_0_70 (.A(A[5]), .ZN(n_0_0_53));
   INV_X1 i_0_0_71 (.A(A[11]), .ZN(n_0_0_54));
   INV_X1 i_0_0_72 (.A(A[15]), .ZN(n_0_0_55));
   INV_X1 i_0_0_73 (.A(B[0]), .ZN(n_0_0_56));
   INV_X1 i_0_0_74 (.A(B[1]), .ZN(n_0_0_57));
   INV_X1 i_0_0_75 (.A(B[3]), .ZN(n_0_0_58));
   INV_X1 i_0_0_76 (.A(B[4]), .ZN(n_0_0_59));
   INV_X1 i_0_0_77 (.A(B[5]), .ZN(n_0_0_60));
   INV_X1 i_0_0_78 (.A(B[11]), .ZN(n_0_0_61));
   INV_X1 i_0_0_79 (.A(B[15]), .ZN(n_0_0_62));
endmodule
