/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Apr 24 23:48:21 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2813677309 */

module datapath(p_0, p_1);
   input [32:0]p_0;
   output [32:0]p_1;

   XOR2_X1 i_0 (.A(p_0[1]), .B(p_0[0]), .Z(p_1[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_1[2]));
   OAI21_X1 i_2 (.A(p_0[2]), .B1(p_0[1]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_0[3]), .B(n_29), .Z(p_1[3]));
   XOR2_X1 i_4 (.A(p_0[4]), .B(n_28), .Z(p_1[4]));
   XOR2_X1 i_5 (.A(p_0[5]), .B(n_27), .Z(p_1[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_1[6]));
   OAI21_X1 i_7 (.A(p_0[6]), .B1(n_27), .B2(p_0[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_0[7]), .B(n_26), .Z(p_1[7]));
   XOR2_X1 i_9 (.A(p_0[8]), .B(n_25), .Z(p_1[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_1[9]));
   OAI21_X1 i_11 (.A(p_0[9]), .B1(n_25), .B2(p_0[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_0[10]), .B(n_24), .Z(p_1[10]));
   XNOR2_X1 i_13 (.A(p_0[11]), .B(n_23), .ZN(p_1[11]));
   XOR2_X1 i_14 (.A(p_0[12]), .B(n_22), .Z(p_1[12]));
   XNOR2_X1 i_15 (.A(p_0[13]), .B(n_21), .ZN(p_1[13]));
   XNOR2_X1 i_16 (.A(p_0[14]), .B(n_20), .ZN(p_1[14]));
   XOR2_X1 i_17 (.A(p_0[15]), .B(n_19), .Z(p_1[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_1[16]));
   OAI21_X1 i_19 (.A(p_0[16]), .B1(n_19), .B2(p_0[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(p_0[17]), .B(n_18), .Z(p_1[17]));
   XOR2_X1 i_21 (.A(p_0[18]), .B(n_17), .Z(p_1[18]));
   XNOR2_X1 i_22 (.A(p_0[19]), .B(n_16), .ZN(p_1[19]));
   XNOR2_X1 i_23 (.A(p_0[20]), .B(n_15), .ZN(p_1[20]));
   XNOR2_X1 i_24 (.A(p_0[21]), .B(n_14), .ZN(p_1[21]));
   XOR2_X1 i_25 (.A(p_0[22]), .B(n_13), .Z(p_1[22]));
   XOR2_X1 i_26 (.A(p_0[23]), .B(n_12), .Z(p_1[23]));
   XNOR2_X1 i_27 (.A(p_0[24]), .B(n_11), .ZN(p_1[24]));
   XNOR2_X1 i_28 (.A(p_0[25]), .B(n_10), .ZN(p_1[25]));
   XOR2_X1 i_29 (.A(p_0[26]), .B(n_9), .Z(p_1[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_1[27]));
   OAI21_X1 i_31 (.A(p_0[27]), .B1(n_9), .B2(p_0[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(p_0[28]), .B(n_8), .Z(p_1[28]));
   XNOR2_X1 i_33 (.A(p_0[29]), .B(n_7), .ZN(p_1[29]));
   XNOR2_X1 i_34 (.A(p_0[30]), .B(n_6), .ZN(p_1[30]));
   XNOR2_X1 i_35 (.A(p_0[31]), .B(n_5), .ZN(p_1[31]));
   NOR2_X1 i_36 (.A1(p_0[31]), .A2(n_5), .ZN(p_1[32]));
   NOR4_X1 i_37 (.A1(n_8), .A2(p_0[28]), .A3(p_0[29]), .A4(p_0[30]), .ZN(n_5));
   NOR3_X1 i_38 (.A1(n_8), .A2(p_0[28]), .A3(p_0[29]), .ZN(n_6));
   NOR2_X1 i_39 (.A1(n_8), .A2(p_0[28]), .ZN(n_7));
   OR3_X1 i_40 (.A1(n_9), .A2(p_0[26]), .A3(p_0[27]), .ZN(n_8));
   NAND2_X1 i_41 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_42 (.A1(n_12), .A2(p_0[23]), .A3(p_0[24]), .ZN(n_10));
   NOR2_X1 i_43 (.A1(n_12), .A2(p_0[23]), .ZN(n_11));
   OR2_X1 i_44 (.A1(n_13), .A2(p_0[22]), .ZN(n_12));
   NAND2_X1 i_45 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_46 (.A1(n_17), .A2(p_0[18]), .A3(p_0[19]), .A4(p_0[20]), .ZN(n_14));
   NOR3_X1 i_47 (.A1(n_17), .A2(p_0[18]), .A3(p_0[19]), .ZN(n_15));
   NOR2_X1 i_48 (.A1(n_17), .A2(p_0[18]), .ZN(n_16));
   OR2_X1 i_49 (.A1(n_18), .A2(p_0[17]), .ZN(n_17));
   OR3_X1 i_50 (.A1(n_19), .A2(p_0[15]), .A3(p_0[16]), .ZN(n_18));
   NAND2_X1 i_51 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_52 (.A1(n_22), .A2(p_0[12]), .A3(p_0[13]), .ZN(n_20));
   NOR2_X1 i_53 (.A1(n_22), .A2(p_0[12]), .ZN(n_21));
   NAND2_X1 i_54 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_55 (.A1(n_24), .A2(p_0[10]), .ZN(n_23));
   OR3_X1 i_56 (.A1(n_25), .A2(p_0[8]), .A3(p_0[9]), .ZN(n_24));
   OR2_X1 i_57 (.A1(n_26), .A2(p_0[7]), .ZN(n_25));
   OR3_X1 i_58 (.A1(n_27), .A2(p_0[5]), .A3(p_0[6]), .ZN(n_26));
   OR2_X1 i_59 (.A1(n_28), .A2(p_0[4]), .ZN(n_27));
   OR2_X1 i_60 (.A1(n_29), .A2(p_0[3]), .ZN(n_28));
   OR3_X1 i_61 (.A1(p_0[2]), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_29));
   INV_X1 i_62 (.A(p_0[11]), .ZN(n_30));
   INV_X1 i_63 (.A(p_0[14]), .ZN(n_31));
   INV_X1 i_64 (.A(p_0[21]), .ZN(n_32));
   INV_X1 i_65 (.A(p_0[25]), .ZN(n_33));
endmodule

module shiftadd(p, a, b, clk, reset);
   output [31:0]p;
   input [15:0]a;
   input [15:0]b;
   input clk;
   input reset;

   wire [15:0]x;
   wire [4:0]i;
   wire n_0_4;
   wire n_0_0;
   wire n_0_5;
   wire n_0_1;
   wire n_0_6;
   wire n_0_2;
   wire n_0_7;
   wire n_0_3;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;

   DFF_X1 \y_reg[32]  (.D(n_87), .CK(n_1), .Q(n_2), .QN());
   DFF_X1 \y_reg[31]  (.D(n_86), .CK(n_1), .Q(p[31]), .QN());
   DFF_X1 \y_reg[30]  (.D(n_85), .CK(n_1), .Q(p[30]), .QN());
   DFF_X1 \y_reg[29]  (.D(n_84), .CK(n_1), .Q(p[29]), .QN());
   DFF_X1 \y_reg[28]  (.D(n_83), .CK(n_1), .Q(p[28]), .QN());
   DFF_X1 \y_reg[27]  (.D(n_82), .CK(n_1), .Q(p[27]), .QN());
   DFF_X1 \y_reg[26]  (.D(n_81), .CK(n_1), .Q(p[26]), .QN());
   DFF_X1 \y_reg[25]  (.D(n_80), .CK(n_1), .Q(p[25]), .QN());
   DFF_X1 \y_reg[24]  (.D(n_79), .CK(n_1), .Q(p[24]), .QN());
   DFF_X1 \y_reg[23]  (.D(n_78), .CK(n_1), .Q(p[23]), .QN());
   DFF_X1 \y_reg[22]  (.D(n_77), .CK(n_1), .Q(p[22]), .QN());
   DFF_X1 \y_reg[21]  (.D(n_76), .CK(n_1), .Q(p[21]), .QN());
   DFF_X1 \y_reg[20]  (.D(n_75), .CK(n_1), .Q(p[20]), .QN());
   DFF_X1 \y_reg[19]  (.D(n_74), .CK(n_1), .Q(p[19]), .QN());
   DFF_X1 \y_reg[18]  (.D(n_73), .CK(n_1), .Q(p[18]), .QN());
   DFF_X1 \y_reg[17]  (.D(n_72), .CK(n_1), .Q(p[17]), .QN());
   DFF_X1 \y_reg[16]  (.D(n_71), .CK(n_1), .Q(p[16]), .QN());
   DFF_X1 \y_reg[15]  (.D(n_70), .CK(n_1), .Q(p[15]), .QN());
   DFF_X1 \y_reg[14]  (.D(n_69), .CK(n_1), .Q(p[14]), .QN());
   DFF_X1 \y_reg[13]  (.D(n_68), .CK(n_1), .Q(p[13]), .QN());
   DFF_X1 \y_reg[12]  (.D(n_67), .CK(n_1), .Q(p[12]), .QN());
   DFF_X1 \y_reg[11]  (.D(n_66), .CK(n_1), .Q(p[11]), .QN());
   DFF_X1 \y_reg[10]  (.D(n_65), .CK(n_1), .Q(p[10]), .QN());
   DFF_X1 \y_reg[9]  (.D(n_64), .CK(n_1), .Q(p[9]), .QN());
   DFF_X1 \y_reg[8]  (.D(n_63), .CK(n_1), .Q(p[8]), .QN());
   DFF_X1 \y_reg[7]  (.D(n_62), .CK(n_1), .Q(p[7]), .QN());
   DFF_X1 \y_reg[6]  (.D(n_61), .CK(n_1), .Q(p[6]), .QN());
   DFF_X1 \y_reg[5]  (.D(n_60), .CK(n_1), .Q(p[5]), .QN());
   DFF_X1 \y_reg[4]  (.D(n_59), .CK(n_1), .Q(p[4]), .QN());
   DFF_X1 \y_reg[3]  (.D(n_58), .CK(n_1), .Q(p[3]), .QN());
   DFF_X1 \y_reg[2]  (.D(n_57), .CK(n_1), .Q(p[2]), .QN());
   DFF_X1 \y_reg[1]  (.D(n_56), .CK(n_1), .Q(p[1]), .QN());
   DFF_X1 \y_reg[0]  (.D(n_55), .CK(n_1), .Q(p[0]), .QN());
   datapath i_4 (.p_0({uc_0, n_119, n_118, n_117, n_116, n_115, n_114, n_113, 
      n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, 
      n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, 
      n_90, n_89, n_88}), .p_1({n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, 
      n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, 
      n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, uc_1}));
   CLKGATETST_X1 clk_gate_x_reg (.CK(clk), .E(reset), .SE(1'b0), .GCK(n_0));
   DFF_X1 \x_reg[15]  (.D(n_54), .CK(n_0), .Q(x[15]), .QN());
   DFF_X1 \x_reg[14]  (.D(n_53), .CK(n_0), .Q(x[14]), .QN());
   DFF_X1 \x_reg[13]  (.D(n_52), .CK(n_0), .Q(x[13]), .QN());
   DFF_X1 \x_reg[12]  (.D(n_51), .CK(n_0), .Q(x[12]), .QN());
   DFF_X1 \x_reg[11]  (.D(n_50), .CK(n_0), .Q(x[11]), .QN());
   DFF_X1 \x_reg[10]  (.D(n_49), .CK(n_0), .Q(x[10]), .QN());
   DFF_X1 \x_reg[9]  (.D(n_48), .CK(n_0), .Q(x[9]), .QN());
   DFF_X1 \x_reg[8]  (.D(n_47), .CK(n_0), .Q(x[8]), .QN());
   DFF_X1 \x_reg[7]  (.D(n_46), .CK(n_0), .Q(x[7]), .QN());
   DFF_X1 \x_reg[6]  (.D(n_45), .CK(n_0), .Q(x[6]), .QN());
   DFF_X1 \x_reg[5]  (.D(n_44), .CK(n_0), .Q(x[5]), .QN());
   DFF_X1 \x_reg[4]  (.D(n_43), .CK(n_0), .Q(x[4]), .QN());
   DFF_X1 \x_reg[3]  (.D(n_42), .CK(n_0), .Q(x[3]), .QN());
   DFF_X1 \x_reg[2]  (.D(n_41), .CK(n_0), .Q(x[2]), .QN());
   DFF_X1 \x_reg[1]  (.D(n_40), .CK(n_0), .Q(x[1]), .QN());
   DFF_X1 \x_reg[0]  (.D(a[0]), .CK(n_0), .Q(x[0]), .QN());
   DFF_X1 \i_reg[4]  (.D(n_39), .CK(n_1), .Q(i[4]), .QN());
   DFF_X1 \i_reg[3]  (.D(n_38), .CK(n_1), .Q(i[3]), .QN());
   DFF_X1 \i_reg[2]  (.D(n_37), .CK(n_1), .Q(i[2]), .QN());
   DFF_X1 \i_reg[1]  (.D(n_36), .CK(n_1), .Q(i[1]), .QN());
   DFF_X1 \i_reg[0]  (.D(n_35), .CK(n_1), .Q(i[0]), .QN());
   CLKGATETST_X1 clk_gate_y_reg (.CK(clk), .E(n_120), .SE(1'b0), .GCK(n_1));
   HA_X1 i_0_0 (.A(i[1]), .B(i[0]), .CO(n_0_0), .S(n_0_4));
   HA_X1 i_0_1 (.A(i[2]), .B(n_0_0), .CO(n_0_1), .S(n_0_5));
   HA_X1 i_0_2 (.A(i[3]), .B(n_0_1), .CO(n_0_2), .S(n_0_6));
   HA_X1 i_0_3 (.A(i[2]), .B(i[1]), .CO(n_0_3), .S(n_0_7));
   HA_X1 i_0_4 (.A(i[3]), .B(n_0_3), .CO(n_0_9), .S(n_0_8));
   AND2_X1 i_0_5 (.A1(n_0_257), .A2(n_0_122), .ZN(n_35));
   NOR2_X1 i_0_6 (.A1(n_0_119), .A2(reset), .ZN(n_36));
   AND2_X1 i_0_7 (.A1(n_0_127), .A2(n_0_257), .ZN(n_37));
   NOR2_X1 i_0_8 (.A1(n_0_117), .A2(reset), .ZN(n_38));
   NOR2_X1 i_0_9 (.A1(reset), .A2(n_0_123), .ZN(n_39));
   XNOR2_X1 i_0_10 (.A(a[1]), .B(n_0_10), .ZN(n_40));
   NAND2_X1 i_0_11 (.A1(a[0]), .A2(n_0_264), .ZN(n_0_10));
   XNOR2_X1 i_0_12 (.A(a[2]), .B(n_0_11), .ZN(n_41));
   OAI21_X1 i_0_13 (.A(n_0_264), .B1(a[0]), .B2(a[1]), .ZN(n_0_11));
   XNOR2_X1 i_0_14 (.A(n_0_253), .B(n_0_12), .ZN(n_42));
   NOR2_X1 i_0_15 (.A1(n_0_34), .A2(n_0_24), .ZN(n_0_12));
   XOR2_X1 i_0_16 (.A(a[4]), .B(n_0_13), .Z(n_43));
   AOI21_X1 i_0_17 (.A(n_0_24), .B1(n_0_34), .B2(n_0_253), .ZN(n_0_13));
   XNOR2_X1 i_0_18 (.A(a[5]), .B(n_0_14), .ZN(n_44));
   NAND2_X1 i_0_19 (.A1(n_0_33), .A2(n_0_264), .ZN(n_0_14));
   XNOR2_X1 i_0_20 (.A(a[6]), .B(n_0_15), .ZN(n_45));
   OAI21_X1 i_0_21 (.A(n_0_264), .B1(n_0_33), .B2(a[5]), .ZN(n_0_15));
   XOR2_X1 i_0_22 (.A(a[7]), .B(n_0_16), .Z(n_46));
   NOR2_X1 i_0_23 (.A1(n_0_32), .A2(n_0_24), .ZN(n_0_16));
   XNOR2_X1 i_0_24 (.A(n_0_255), .B(n_0_17), .ZN(n_47));
   NOR2_X1 i_0_25 (.A1(n_0_31), .A2(n_0_24), .ZN(n_0_17));
   XNOR2_X1 i_0_26 (.A(a[9]), .B(n_0_18), .ZN(n_48));
   NAND2_X1 i_0_27 (.A1(n_0_30), .A2(n_0_264), .ZN(n_0_18));
   XNOR2_X1 i_0_28 (.A(a[10]), .B(n_0_19), .ZN(n_49));
   NAND2_X1 i_0_29 (.A1(n_0_29), .A2(n_0_264), .ZN(n_0_19));
   XNOR2_X1 i_0_30 (.A(a[11]), .B(n_0_20), .ZN(n_50));
   NAND2_X1 i_0_31 (.A1(n_0_28), .A2(n_0_264), .ZN(n_0_20));
   XNOR2_X1 i_0_32 (.A(a[12]), .B(n_0_21), .ZN(n_51));
   OAI21_X1 i_0_33 (.A(n_0_264), .B1(n_0_28), .B2(a[11]), .ZN(n_0_21));
   XNOR2_X1 i_0_34 (.A(n_0_256), .B(n_0_22), .ZN(n_52));
   NOR2_X1 i_0_35 (.A1(n_0_27), .A2(n_0_24), .ZN(n_0_22));
   XOR2_X1 i_0_36 (.A(a[14]), .B(n_0_23), .Z(n_53));
   AOI21_X1 i_0_37 (.A(n_0_24), .B1(n_0_27), .B2(n_0_256), .ZN(n_0_23));
   NAND2_X1 i_0_38 (.A1(reset), .A2(a[15]), .ZN(n_0_24));
   AND2_X1 i_0_39 (.A1(n_0_25), .A2(a[15]), .ZN(n_54));
   OAI21_X1 i_0_40 (.A(reset), .B1(n_0_26), .B2(a[14]), .ZN(n_0_25));
   NAND2_X1 i_0_41 (.A1(n_0_27), .A2(n_0_256), .ZN(n_0_26));
   NOR3_X1 i_0_42 (.A1(n_0_28), .A2(a[11]), .A3(a[12]), .ZN(n_0_27));
   OR2_X1 i_0_43 (.A1(n_0_29), .A2(a[10]), .ZN(n_0_28));
   OR2_X1 i_0_44 (.A1(n_0_30), .A2(a[9]), .ZN(n_0_29));
   NAND2_X1 i_0_45 (.A1(n_0_31), .A2(n_0_255), .ZN(n_0_30));
   NOR4_X1 i_0_46 (.A1(n_0_33), .A2(a[5]), .A3(a[6]), .A4(a[7]), .ZN(n_0_31));
   NOR3_X1 i_0_47 (.A1(n_0_33), .A2(a[5]), .A3(a[6]), .ZN(n_0_32));
   NAND3_X1 i_0_48 (.A1(n_0_34), .A2(n_0_253), .A3(n_0_254), .ZN(n_0_33));
   NOR3_X1 i_0_49 (.A1(a[2]), .A2(a[1]), .A3(a[0]), .ZN(n_0_34));
   INV_X1 i_0_50 (.A(n_0_35), .ZN(n_55));
   AOI22_X1 i_0_51 (.A1(n_88), .A2(n_0_115), .B1(b[0]), .B2(reset), .ZN(n_0_35));
   OAI21_X1 i_0_52 (.A(n_0_36), .B1(n_0_37), .B2(n_0_257), .ZN(n_56));
   AOI22_X1 i_0_53 (.A1(n_89), .A2(n_0_114), .B1(n_0_112), .B2(n_3), .ZN(n_0_36));
   XOR2_X1 i_0_54 (.A(b[1]), .B(n_0_38), .Z(n_0_37));
   NAND2_X1 i_0_55 (.A1(b[15]), .A2(b[0]), .ZN(n_0_38));
   INV_X1 i_0_56 (.A(n_0_39), .ZN(n_57));
   AOI222_X1 i_0_57 (.A1(n_90), .A2(n_0_114), .B1(n_0_112), .B2(n_4), .C1(reset), 
      .C2(n_0_40), .ZN(n_0_39));
   XNOR2_X1 i_0_58 (.A(b[2]), .B(n_0_41), .ZN(n_0_40));
   OAI21_X1 i_0_59 (.A(b[15]), .B1(b[1]), .B2(b[0]), .ZN(n_0_41));
   OAI21_X1 i_0_60 (.A(n_0_42), .B1(n_0_43), .B2(n_0_44), .ZN(n_58));
   AOI22_X1 i_0_61 (.A1(n_91), .A2(n_0_114), .B1(n_0_112), .B2(n_5), .ZN(n_0_42));
   NAND2_X1 i_0_62 (.A1(n_0_45), .A2(reset), .ZN(n_0_43));
   AOI21_X1 i_0_63 (.A(b[3]), .B1(n_0_93), .B2(b[15]), .ZN(n_0_44));
   NAND3_X1 i_0_64 (.A1(n_0_93), .A2(b[3]), .A3(b[15]), .ZN(n_0_45));
   OAI21_X1 i_0_65 (.A(n_0_46), .B1(n_0_47), .B2(n_0_257), .ZN(n_59));
   AOI22_X1 i_0_66 (.A1(n_92), .A2(n_0_114), .B1(n_0_112), .B2(n_6), .ZN(n_0_46));
   INV_X1 i_0_67 (.A(n_0_48), .ZN(n_0_47));
   XNOR2_X1 i_0_68 (.A(b[4]), .B(n_0_49), .ZN(n_0_48));
   OAI21_X1 i_0_69 (.A(b[15]), .B1(n_0_93), .B2(b[3]), .ZN(n_0_49));
   OAI21_X1 i_0_70 (.A(n_0_50), .B1(n_0_51), .B2(n_0_52), .ZN(n_60));
   AOI22_X1 i_0_71 (.A1(n_93), .A2(n_0_114), .B1(n_0_112), .B2(n_7), .ZN(n_0_50));
   NAND2_X1 i_0_72 (.A1(n_0_53), .A2(reset), .ZN(n_0_51));
   AOI21_X1 i_0_73 (.A(b[5]), .B1(n_0_92), .B2(b[15]), .ZN(n_0_52));
   NAND3_X1 i_0_74 (.A1(n_0_92), .A2(b[5]), .A3(b[15]), .ZN(n_0_53));
   OAI21_X1 i_0_75 (.A(n_0_54), .B1(n_0_55), .B2(n_0_257), .ZN(n_61));
   AOI22_X1 i_0_76 (.A1(n_94), .A2(n_0_114), .B1(n_0_112), .B2(n_8), .ZN(n_0_54));
   INV_X1 i_0_77 (.A(n_0_56), .ZN(n_0_55));
   XNOR2_X1 i_0_78 (.A(b[6]), .B(n_0_57), .ZN(n_0_56));
   OAI21_X1 i_0_79 (.A(b[15]), .B1(n_0_92), .B2(b[5]), .ZN(n_0_57));
   INV_X1 i_0_80 (.A(n_0_58), .ZN(n_62));
   AOI222_X1 i_0_81 (.A1(n_95), .A2(n_0_114), .B1(n_0_112), .B2(n_9), .C1(reset), 
      .C2(n_0_59), .ZN(n_0_58));
   XNOR2_X1 i_0_82 (.A(b[7]), .B(n_0_60), .ZN(n_0_59));
   NAND2_X1 i_0_83 (.A1(n_0_91), .A2(b[15]), .ZN(n_0_60));
   INV_X1 i_0_84 (.A(n_0_61), .ZN(n_63));
   AOI222_X1 i_0_85 (.A1(n_96), .A2(n_0_114), .B1(n_0_112), .B2(n_10), .C1(reset), 
      .C2(n_0_62), .ZN(n_0_61));
   XNOR2_X1 i_0_86 (.A(n_0_260), .B(n_0_63), .ZN(n_0_62));
   NOR2_X1 i_0_87 (.A1(n_0_90), .A2(n_0_261), .ZN(n_0_63));
   INV_X1 i_0_88 (.A(n_0_64), .ZN(n_64));
   AOI222_X1 i_0_89 (.A1(n_97), .A2(n_0_114), .B1(n_0_112), .B2(n_11), .C1(reset), 
      .C2(n_0_65), .ZN(n_0_64));
   XNOR2_X1 i_0_90 (.A(b[9]), .B(n_0_66), .ZN(n_0_65));
   NAND2_X1 i_0_91 (.A1(n_0_89), .A2(b[15]), .ZN(n_0_66));
   INV_X1 i_0_92 (.A(n_0_67), .ZN(n_65));
   AOI222_X1 i_0_93 (.A1(n_98), .A2(n_0_114), .B1(n_0_112), .B2(n_12), .C1(reset), 
      .C2(n_0_68), .ZN(n_0_67));
   XNOR2_X1 i_0_94 (.A(b[10]), .B(n_0_69), .ZN(n_0_68));
   NAND2_X1 i_0_95 (.A1(n_0_88), .A2(b[15]), .ZN(n_0_69));
   INV_X1 i_0_96 (.A(n_0_70), .ZN(n_66));
   AOI222_X1 i_0_97 (.A1(n_99), .A2(n_0_114), .B1(n_0_112), .B2(n_13), .C1(reset), 
      .C2(n_0_71), .ZN(n_0_70));
   XNOR2_X1 i_0_98 (.A(b[11]), .B(n_0_72), .ZN(n_0_71));
   NAND2_X1 i_0_99 (.A1(n_0_87), .A2(b[15]), .ZN(n_0_72));
   INV_X1 i_0_100 (.A(n_0_73), .ZN(n_67));
   AOI222_X1 i_0_101 (.A1(n_100), .A2(n_0_114), .B1(n_0_112), .B2(n_14), 
      .C1(reset), .C2(n_0_74), .ZN(n_0_73));
   XNOR2_X1 i_0_102 (.A(b[12]), .B(n_0_75), .ZN(n_0_74));
   NAND2_X1 i_0_103 (.A1(n_0_86), .A2(b[15]), .ZN(n_0_75));
   INV_X1 i_0_104 (.A(n_0_76), .ZN(n_68));
   AOI222_X1 i_0_105 (.A1(n_101), .A2(n_0_114), .B1(n_0_112), .B2(n_15), 
      .C1(reset), .C2(n_0_77), .ZN(n_0_76));
   XNOR2_X1 i_0_106 (.A(b[13]), .B(n_0_78), .ZN(n_0_77));
   NAND2_X1 i_0_107 (.A1(n_0_85), .A2(b[15]), .ZN(n_0_78));
   NAND2_X1 i_0_108 (.A1(n_0_79), .A2(n_0_81), .ZN(n_69));
   AOI22_X1 i_0_109 (.A1(reset), .A2(n_0_80), .B1(n_0_114), .B2(n_102), .ZN(
      n_0_79));
   XNOR2_X1 i_0_110 (.A(b[14]), .B(n_0_82), .ZN(n_0_80));
   NAND2_X1 i_0_111 (.A1(n_16), .A2(n_0_112), .ZN(n_0_81));
   NAND2_X1 i_0_112 (.A1(n_0_84), .A2(b[15]), .ZN(n_0_82));
   OAI21_X1 i_0_113 (.A(n_0_94), .B1(n_0_84), .B2(n_0_83), .ZN(n_70));
   OR3_X1 i_0_114 (.A1(n_0_261), .A2(n_0_257), .A3(b[14]), .ZN(n_0_83));
   OR2_X1 i_0_115 (.A1(n_0_85), .A2(b[13]), .ZN(n_0_84));
   OR2_X1 i_0_116 (.A1(n_0_86), .A2(b[12]), .ZN(n_0_85));
   OR2_X1 i_0_117 (.A1(n_0_87), .A2(b[11]), .ZN(n_0_86));
   OR2_X1 i_0_118 (.A1(n_0_88), .A2(b[10]), .ZN(n_0_87));
   OR2_X1 i_0_119 (.A1(n_0_89), .A2(b[9]), .ZN(n_0_88));
   NAND2_X1 i_0_120 (.A1(n_0_90), .A2(n_0_260), .ZN(n_0_89));
   NOR2_X1 i_0_121 (.A1(n_0_91), .A2(b[7]), .ZN(n_0_90));
   OR3_X1 i_0_122 (.A1(n_0_92), .A2(b[5]), .A3(b[6]), .ZN(n_0_91));
   OR3_X1 i_0_123 (.A1(n_0_93), .A2(b[3]), .A3(b[4]), .ZN(n_0_92));
   OR3_X1 i_0_124 (.A1(b[2]), .A2(b[1]), .A3(b[0]), .ZN(n_0_93));
   AOI22_X1 i_0_125 (.A1(n_0_114), .A2(n_103), .B1(n_17), .B2(n_0_112), .ZN(
      n_0_94));
   INV_X1 i_0_126 (.A(n_0_95), .ZN(n_71));
   AOI22_X1 i_0_127 (.A1(n_0_114), .A2(n_104), .B1(n_18), .B2(n_0_112), .ZN(
      n_0_95));
   INV_X1 i_0_128 (.A(n_0_96), .ZN(n_72));
   AOI22_X1 i_0_129 (.A1(n_0_114), .A2(n_105), .B1(n_19), .B2(n_0_112), .ZN(
      n_0_96));
   INV_X1 i_0_130 (.A(n_0_97), .ZN(n_73));
   AOI22_X1 i_0_131 (.A1(n_106), .A2(n_0_114), .B1(n_0_112), .B2(n_20), .ZN(
      n_0_97));
   INV_X1 i_0_132 (.A(n_0_98), .ZN(n_74));
   AOI22_X1 i_0_133 (.A1(n_107), .A2(n_0_114), .B1(n_0_112), .B2(n_21), .ZN(
      n_0_98));
   INV_X1 i_0_134 (.A(n_0_99), .ZN(n_75));
   AOI22_X1 i_0_135 (.A1(n_108), .A2(n_0_114), .B1(n_0_112), .B2(n_22), .ZN(
      n_0_99));
   INV_X1 i_0_136 (.A(n_0_100), .ZN(n_76));
   AOI22_X1 i_0_137 (.A1(n_109), .A2(n_0_114), .B1(n_0_112), .B2(n_23), .ZN(
      n_0_100));
   INV_X1 i_0_138 (.A(n_0_101), .ZN(n_77));
   AOI22_X1 i_0_139 (.A1(n_110), .A2(n_0_114), .B1(n_0_112), .B2(n_24), .ZN(
      n_0_101));
   INV_X1 i_0_140 (.A(n_0_102), .ZN(n_78));
   AOI22_X1 i_0_141 (.A1(n_111), .A2(n_0_114), .B1(n_0_112), .B2(n_25), .ZN(
      n_0_102));
   INV_X1 i_0_142 (.A(n_0_103), .ZN(n_79));
   AOI22_X1 i_0_143 (.A1(n_112), .A2(n_0_114), .B1(n_0_112), .B2(n_26), .ZN(
      n_0_103));
   INV_X1 i_0_144 (.A(n_0_104), .ZN(n_80));
   AOI22_X1 i_0_145 (.A1(n_113), .A2(n_0_114), .B1(n_0_112), .B2(n_27), .ZN(
      n_0_104));
   INV_X1 i_0_146 (.A(n_0_105), .ZN(n_81));
   AOI22_X1 i_0_147 (.A1(n_114), .A2(n_0_114), .B1(n_0_112), .B2(n_28), .ZN(
      n_0_105));
   INV_X1 i_0_148 (.A(n_0_106), .ZN(n_82));
   AOI22_X1 i_0_149 (.A1(n_115), .A2(n_0_114), .B1(n_0_112), .B2(n_29), .ZN(
      n_0_106));
   INV_X1 i_0_150 (.A(n_0_107), .ZN(n_83));
   AOI22_X1 i_0_151 (.A1(n_116), .A2(n_0_114), .B1(n_0_112), .B2(n_30), .ZN(
      n_0_107));
   INV_X1 i_0_152 (.A(n_0_108), .ZN(n_84));
   AOI22_X1 i_0_153 (.A1(n_117), .A2(n_0_114), .B1(n_0_112), .B2(n_31), .ZN(
      n_0_108));
   INV_X1 i_0_154 (.A(n_0_109), .ZN(n_85));
   AOI22_X1 i_0_155 (.A1(n_118), .A2(n_0_114), .B1(n_0_112), .B2(n_32), .ZN(
      n_0_109));
   NAND2_X1 i_0_156 (.A1(n_0_113), .A2(n_0_110), .ZN(n_86));
   NAND2_X1 i_0_157 (.A1(n_33), .A2(n_0_112), .ZN(n_0_110));
   NAND2_X1 i_0_158 (.A1(n_0_113), .A2(n_0_111), .ZN(n_87));
   NAND2_X1 i_0_159 (.A1(n_34), .A2(n_0_112), .ZN(n_0_111));
   NOR2_X1 i_0_160 (.A1(n_0_116), .A2(reset), .ZN(n_0_112));
   NAND2_X1 i_0_161 (.A1(n_119), .A2(n_0_114), .ZN(n_0_113));
   AND2_X1 i_0_162 (.A1(n_0_116), .A2(n_0_115), .ZN(n_0_114));
   NOR2_X1 i_0_163 (.A1(i[4]), .A2(reset), .ZN(n_0_115));
   NAND4_X1 i_0_164 (.A1(n_0_126), .A2(n_0_121), .A3(n_0_119), .A4(n_0_117), 
      .ZN(n_0_116));
   OAI21_X1 i_0_165 (.A(n_0_118), .B1(n_0_194), .B2(n_0_8), .ZN(n_0_117));
   OR2_X1 i_0_166 (.A1(n_0_6), .A2(n_0_262), .ZN(n_0_118));
   OAI21_X1 i_0_167 (.A(n_0_120), .B1(n_0_262), .B2(n_0_4), .ZN(n_0_119));
   NAND2_X1 i_0_168 (.A1(i[1]), .A2(n_0_262), .ZN(n_0_120));
   NOR2_X1 i_0_169 (.A1(n_0_123), .A2(n_0_122), .ZN(n_0_121));
   XNOR2_X1 i_0_170 (.A(i[0]), .B(n_0_262), .ZN(n_0_122));
   AOI21_X1 i_0_171 (.A(n_0_124), .B1(n_0_262), .B2(n_0_9), .ZN(n_0_123));
   NOR2_X1 i_0_172 (.A1(n_0_262), .A2(n_0_125), .ZN(n_0_124));
   XNOR2_X1 i_0_173 (.A(i[4]), .B(n_0_2), .ZN(n_0_125));
   AOI211_X1 i_0_174 (.A(n_0_128), .B(n_0_127), .C1(b[15]), .C2(a[15]), .ZN(
      n_0_126));
   MUX2_X1 i_0_175 (.A(n_0_5), .B(n_0_7), .S(n_0_262), .Z(n_0_127));
   OAI21_X1 i_0_176 (.A(n_0_259), .B1(a[15]), .B2(b[15]), .ZN(n_0_128));
   INV_X1 i_0_177 (.A(n_0_129), .ZN(n_88));
   AOI21_X1 i_0_178 (.A(p[1]), .B1(n_0_195), .B2(p[2]), .ZN(n_0_129));
   MUX2_X1 i_0_179 (.A(p[2]), .B(p[3]), .S(n_0_262), .Z(n_89));
   MUX2_X1 i_0_180 (.A(p[3]), .B(p[4]), .S(n_0_262), .Z(n_90));
   MUX2_X1 i_0_181 (.A(p[4]), .B(p[5]), .S(n_0_262), .Z(n_91));
   MUX2_X1 i_0_182 (.A(p[5]), .B(p[6]), .S(n_0_262), .Z(n_92));
   MUX2_X1 i_0_183 (.A(p[6]), .B(p[7]), .S(n_0_262), .Z(n_93));
   MUX2_X1 i_0_184 (.A(p[7]), .B(p[8]), .S(n_0_262), .Z(n_94));
   MUX2_X1 i_0_185 (.A(p[8]), .B(p[9]), .S(n_0_262), .Z(n_95));
   MUX2_X1 i_0_186 (.A(p[9]), .B(p[10]), .S(n_0_262), .Z(n_96));
   MUX2_X1 i_0_187 (.A(p[10]), .B(p[11]), .S(n_0_262), .Z(n_97));
   MUX2_X1 i_0_188 (.A(p[11]), .B(p[12]), .S(n_0_262), .Z(n_98));
   MUX2_X1 i_0_189 (.A(p[12]), .B(p[13]), .S(n_0_262), .Z(n_99));
   MUX2_X1 i_0_190 (.A(p[13]), .B(p[14]), .S(n_0_262), .Z(n_100));
   MUX2_X1 i_0_191 (.A(p[14]), .B(p[15]), .S(n_0_262), .Z(n_101));
   OAI21_X1 i_0_192 (.A(n_0_130), .B1(n_0_133), .B2(n_0_193), .ZN(n_102));
   AOI22_X1 i_0_193 (.A1(p[16]), .A2(n_0_191), .B1(n_0_194), .B2(p[15]), 
      .ZN(n_0_130));
   INV_X1 i_0_194 (.A(n_0_131), .ZN(n_103));
   AOI221_X1 i_0_195 (.A(n_0_132), .B1(n_0_192), .B2(p[16]), .C1(p[17]), 
      .C2(n_0_191), .ZN(n_0_131));
   OAI22_X1 i_0_196 (.A1(n_0_193), .A2(n_0_134), .B1(n_0_133), .B2(n_0_189), 
      .ZN(n_0_132));
   XNOR2_X1 i_0_197 (.A(p[16]), .B(x[0]), .ZN(n_0_133));
   OAI211_X1 i_0_198 (.A(n_0_136), .B(n_0_135), .C1(n_0_134), .C2(n_0_189), 
      .ZN(n_104));
   XNOR2_X1 i_0_199 (.A(n_0_236), .B(n_0_235), .ZN(n_0_134));
   AOI22_X1 i_0_200 (.A1(p[17]), .A2(n_0_192), .B1(n_0_191), .B2(p[18]), 
      .ZN(n_0_135));
   NAND2_X1 i_0_201 (.A1(n_0_138), .A2(n_0_263), .ZN(n_0_136));
   OAI211_X1 i_0_202 (.A(n_0_137), .B(n_0_140), .C1(n_0_143), .C2(n_0_193), 
      .ZN(n_105));
   NAND3_X1 i_0_203 (.A1(n_0_138), .A2(p[0]), .A3(n_0_194), .ZN(n_0_137));
   XNOR2_X1 i_0_204 (.A(n_0_234), .B(n_0_139), .ZN(n_0_138));
   XNOR2_X1 i_0_205 (.A(p[18]), .B(x[2]), .ZN(n_0_139));
   AOI22_X1 i_0_206 (.A1(p[18]), .A2(n_0_192), .B1(n_0_191), .B2(p[19]), 
      .ZN(n_0_140));
   OAI21_X1 i_0_207 (.A(n_0_141), .B1(n_0_147), .B2(n_0_193), .ZN(n_106));
   AOI221_X1 i_0_208 (.A(n_0_142), .B1(n_0_192), .B2(p[19]), .C1(p[20]), 
      .C2(n_0_191), .ZN(n_0_141));
   NOR2_X1 i_0_209 (.A1(n_0_143), .A2(n_0_189), .ZN(n_0_142));
   XNOR2_X1 i_0_210 (.A(n_0_231), .B(n_0_144), .ZN(n_0_143));
   XOR2_X1 i_0_211 (.A(p[19]), .B(x[3]), .Z(n_0_144));
   OAI21_X1 i_0_212 (.A(n_0_145), .B1(n_0_151), .B2(n_0_193), .ZN(n_107));
   AOI221_X1 i_0_213 (.A(n_0_146), .B1(n_0_192), .B2(p[20]), .C1(p[21]), 
      .C2(n_0_191), .ZN(n_0_145));
   NOR2_X1 i_0_214 (.A1(n_0_189), .A2(n_0_147), .ZN(n_0_146));
   XOR2_X1 i_0_215 (.A(x[4]), .B(n_0_148), .Z(n_0_147));
   NAND2_X1 i_0_216 (.A1(n_0_226), .A2(n_0_225), .ZN(n_0_148));
   OAI21_X1 i_0_217 (.A(n_0_149), .B1(n_0_155), .B2(n_0_193), .ZN(n_108));
   AOI221_X1 i_0_218 (.A(n_0_150), .B1(n_0_192), .B2(p[21]), .C1(p[22]), 
      .C2(n_0_191), .ZN(n_0_149));
   NOR2_X1 i_0_219 (.A1(n_0_189), .A2(n_0_151), .ZN(n_0_150));
   XNOR2_X1 i_0_220 (.A(n_0_224), .B(n_0_152), .ZN(n_0_151));
   OR2_X1 i_0_221 (.A1(n_0_240), .A2(n_0_238), .ZN(n_0_152));
   OAI21_X1 i_0_222 (.A(n_0_153), .B1(n_0_157), .B2(n_0_193), .ZN(n_109));
   AOI221_X1 i_0_223 (.A(n_0_154), .B1(n_0_192), .B2(p[22]), .C1(p[23]), 
      .C2(n_0_191), .ZN(n_0_153));
   NOR2_X1 i_0_224 (.A1(n_0_189), .A2(n_0_155), .ZN(n_0_154));
   XNOR2_X1 i_0_225 (.A(n_0_223), .B(n_0_156), .ZN(n_0_155));
   XOR2_X1 i_0_226 (.A(p[22]), .B(x[6]), .Z(n_0_156));
   OAI211_X1 i_0_227 (.A(n_0_160), .B(n_0_159), .C1(n_0_157), .C2(n_0_189), 
      .ZN(n_110));
   XNOR2_X1 i_0_228 (.A(n_0_220), .B(n_0_158), .ZN(n_0_157));
   OR2_X1 i_0_229 (.A1(n_0_243), .A2(n_0_241), .ZN(n_0_158));
   AOI22_X1 i_0_230 (.A1(p[23]), .A2(n_0_192), .B1(n_0_191), .B2(p[24]), 
      .ZN(n_0_159));
   NAND2_X1 i_0_231 (.A1(n_0_263), .A2(n_0_162), .ZN(n_0_160));
   OAI211_X1 i_0_232 (.A(n_0_161), .B(n_0_164), .C1(n_0_167), .C2(n_0_193), 
      .ZN(n_111));
   NAND3_X1 i_0_233 (.A1(p[0]), .A2(n_0_162), .A3(n_0_194), .ZN(n_0_161));
   XNOR2_X1 i_0_234 (.A(n_0_219), .B(n_0_163), .ZN(n_0_162));
   XNOR2_X1 i_0_235 (.A(p[24]), .B(x[8]), .ZN(n_0_163));
   AOI22_X1 i_0_236 (.A1(p[24]), .A2(n_0_192), .B1(n_0_191), .B2(p[25]), 
      .ZN(n_0_164));
   OAI21_X1 i_0_237 (.A(n_0_165), .B1(n_0_171), .B2(n_0_193), .ZN(n_112));
   AOI221_X1 i_0_238 (.A(n_0_166), .B1(n_0_192), .B2(p[25]), .C1(p[26]), 
      .C2(n_0_191), .ZN(n_0_165));
   NOR2_X1 i_0_239 (.A1(n_0_189), .A2(n_0_167), .ZN(n_0_166));
   XNOR2_X1 i_0_240 (.A(n_0_216), .B(n_0_168), .ZN(n_0_167));
   OR2_X1 i_0_241 (.A1(n_0_246), .A2(n_0_244), .ZN(n_0_168));
   OAI21_X1 i_0_242 (.A(n_0_169), .B1(n_0_173), .B2(n_0_193), .ZN(n_113));
   AOI221_X1 i_0_243 (.A(n_0_170), .B1(n_0_192), .B2(p[26]), .C1(p[27]), 
      .C2(n_0_191), .ZN(n_0_169));
   NOR2_X1 i_0_244 (.A1(n_0_189), .A2(n_0_171), .ZN(n_0_170));
   XNOR2_X1 i_0_245 (.A(n_0_215), .B(n_0_172), .ZN(n_0_171));
   XOR2_X1 i_0_246 (.A(p[26]), .B(x[10]), .Z(n_0_172));
   OAI211_X1 i_0_247 (.A(n_0_176), .B(n_0_175), .C1(n_0_173), .C2(n_0_189), 
      .ZN(n_114));
   XNOR2_X1 i_0_248 (.A(n_0_212), .B(n_0_174), .ZN(n_0_173));
   OR2_X1 i_0_249 (.A1(n_0_249), .A2(n_0_247), .ZN(n_0_174));
   AOI22_X1 i_0_250 (.A1(p[27]), .A2(n_0_192), .B1(n_0_191), .B2(p[28]), 
      .ZN(n_0_175));
   NAND2_X1 i_0_251 (.A1(n_0_263), .A2(n_0_178), .ZN(n_0_176));
   OAI211_X1 i_0_252 (.A(n_0_177), .B(n_0_180), .C1(n_0_183), .C2(n_0_193), 
      .ZN(n_115));
   NAND3_X1 i_0_253 (.A1(p[0]), .A2(n_0_178), .A3(n_0_194), .ZN(n_0_177));
   XNOR2_X1 i_0_254 (.A(n_0_211), .B(n_0_179), .ZN(n_0_178));
   XNOR2_X1 i_0_255 (.A(p[28]), .B(x[12]), .ZN(n_0_179));
   AOI22_X1 i_0_256 (.A1(p[28]), .A2(n_0_192), .B1(n_0_191), .B2(p[29]), 
      .ZN(n_0_180));
   OAI21_X1 i_0_257 (.A(n_0_181), .B1(n_0_187), .B2(n_0_193), .ZN(n_116));
   AOI221_X1 i_0_258 (.A(n_0_182), .B1(n_0_192), .B2(p[29]), .C1(p[30]), 
      .C2(n_0_191), .ZN(n_0_181));
   NOR2_X1 i_0_259 (.A1(n_0_189), .A2(n_0_183), .ZN(n_0_182));
   XNOR2_X1 i_0_260 (.A(n_0_208), .B(n_0_184), .ZN(n_0_183));
   OR2_X1 i_0_261 (.A1(n_0_252), .A2(n_0_250), .ZN(n_0_184));
   OAI21_X1 i_0_262 (.A(n_0_185), .B1(n_0_193), .B2(n_0_200), .ZN(n_117));
   AOI221_X1 i_0_263 (.A(n_0_186), .B1(n_0_192), .B2(p[30]), .C1(p[31]), 
      .C2(n_0_191), .ZN(n_0_185));
   NOR2_X1 i_0_264 (.A1(n_0_189), .A2(n_0_187), .ZN(n_0_186));
   XNOR2_X1 i_0_265 (.A(n_0_207), .B(n_0_188), .ZN(n_0_187));
   XOR2_X1 i_0_266 (.A(p[30]), .B(x[14]), .Z(n_0_188));
   OAI221_X1 i_0_267 (.A(n_0_190), .B1(n_0_189), .B2(n_0_200), .C1(n_0_199), 
      .C2(n_0_193), .ZN(n_118));
   NAND2_X1 i_0_268 (.A1(n_0_194), .A2(p[0]), .ZN(n_0_189));
   AOI22_X1 i_0_269 (.A1(p[31]), .A2(n_0_192), .B1(n_0_191), .B2(n_2), .ZN(
      n_0_190));
   NOR2_X1 i_0_270 (.A1(n_0_194), .A2(p[0]), .ZN(n_0_191));
   NOR2_X1 i_0_271 (.A1(p[0]), .A2(n_0_262), .ZN(n_0_192));
   NAND2_X1 i_0_272 (.A1(p[0]), .A2(n_0_262), .ZN(n_0_193));
   OR2_X1 i_0_273 (.A1(n_0_196), .A2(p[1]), .ZN(n_0_194));
   INV_X1 i_0_274 (.A(n_0_196), .ZN(n_0_195));
   NAND2_X1 i_0_275 (.A1(n_0_259), .A2(n_0_197), .ZN(n_0_196));
   NAND4_X1 i_0_276 (.A1(i[3]), .A2(i[2]), .A3(i[1]), .A4(i[0]), .ZN(n_0_197));
   AOI21_X1 i_0_277 (.A(n_0_198), .B1(n_0_199), .B2(p[0]), .ZN(n_119));
   NOR2_X1 i_0_278 (.A1(n_2), .A2(p[0]), .ZN(n_0_198));
   MUX2_X1 i_0_279 (.A(n_0_203), .B(n_0_202), .S(n_0_204), .Z(n_0_199));
   XNOR2_X1 i_0_280 (.A(n_0_204), .B(n_0_201), .ZN(n_0_200));
   NAND2_X1 i_0_281 (.A1(n_0_203), .A2(n_0_202), .ZN(n_0_201));
   NAND2_X1 i_0_282 (.A1(p[31]), .A2(x[15]), .ZN(n_0_202));
   OR2_X1 i_0_283 (.A1(p[31]), .A2(x[15]), .ZN(n_0_203));
   OAI21_X1 i_0_284 (.A(n_0_205), .B1(n_0_207), .B2(p[30]), .ZN(n_0_204));
   INV_X1 i_0_285 (.A(n_0_206), .ZN(n_0_205));
   AOI21_X1 i_0_286 (.A(x[14]), .B1(n_0_207), .B2(p[30]), .ZN(n_0_206));
   OAI21_X1 i_0_287 (.A(n_0_251), .B1(n_0_208), .B2(n_0_252), .ZN(n_0_207));
   OAI21_X1 i_0_288 (.A(n_0_209), .B1(n_0_211), .B2(p[28]), .ZN(n_0_208));
   INV_X1 i_0_289 (.A(n_0_210), .ZN(n_0_209));
   AOI21_X1 i_0_290 (.A(x[12]), .B1(n_0_211), .B2(p[28]), .ZN(n_0_210));
   OAI21_X1 i_0_291 (.A(n_0_248), .B1(n_0_212), .B2(n_0_249), .ZN(n_0_211));
   OAI21_X1 i_0_292 (.A(n_0_213), .B1(n_0_215), .B2(p[26]), .ZN(n_0_212));
   INV_X1 i_0_293 (.A(n_0_214), .ZN(n_0_213));
   AOI21_X1 i_0_294 (.A(x[10]), .B1(n_0_215), .B2(p[26]), .ZN(n_0_214));
   OAI21_X1 i_0_295 (.A(n_0_245), .B1(n_0_216), .B2(n_0_246), .ZN(n_0_215));
   OAI21_X1 i_0_296 (.A(n_0_217), .B1(n_0_219), .B2(p[24]), .ZN(n_0_216));
   INV_X1 i_0_297 (.A(n_0_218), .ZN(n_0_217));
   AOI21_X1 i_0_298 (.A(x[8]), .B1(n_0_219), .B2(p[24]), .ZN(n_0_218));
   OAI21_X1 i_0_299 (.A(n_0_242), .B1(n_0_220), .B2(n_0_243), .ZN(n_0_219));
   OAI21_X1 i_0_300 (.A(n_0_221), .B1(n_0_223), .B2(p[22]), .ZN(n_0_220));
   INV_X1 i_0_301 (.A(n_0_222), .ZN(n_0_221));
   AOI21_X1 i_0_302 (.A(x[6]), .B1(n_0_223), .B2(p[22]), .ZN(n_0_222));
   OAI21_X1 i_0_303 (.A(n_0_239), .B1(n_0_224), .B2(n_0_240), .ZN(n_0_223));
   OAI21_X1 i_0_304 (.A(n_0_225), .B1(n_0_227), .B2(x[4]), .ZN(n_0_224));
   NAND2_X1 i_0_305 (.A1(n_0_258), .A2(n_0_228), .ZN(n_0_225));
   INV_X1 i_0_306 (.A(n_0_227), .ZN(n_0_226));
   NOR2_X1 i_0_307 (.A1(n_0_258), .A2(n_0_228), .ZN(n_0_227));
   OAI21_X1 i_0_308 (.A(n_0_229), .B1(x[3]), .B2(p[19]), .ZN(n_0_228));
   INV_X1 i_0_309 (.A(n_0_230), .ZN(n_0_229));
   AOI21_X1 i_0_310 (.A(n_0_231), .B1(x[3]), .B2(p[19]), .ZN(n_0_230));
   NOR2_X1 i_0_311 (.A1(n_0_233), .A2(n_0_232), .ZN(n_0_231));
   NOR2_X1 i_0_312 (.A1(n_0_234), .A2(p[18]), .ZN(n_0_232));
   AOI21_X1 i_0_313 (.A(x[2]), .B1(n_0_234), .B2(p[18]), .ZN(n_0_233));
   OAI21_X1 i_0_314 (.A(n_0_237), .B1(n_0_236), .B2(n_0_235), .ZN(n_0_234));
   XNOR2_X1 i_0_315 (.A(p[17]), .B(x[1]), .ZN(n_0_235));
   NAND2_X1 i_0_316 (.A1(p[16]), .A2(x[0]), .ZN(n_0_236));
   NAND2_X1 i_0_317 (.A1(p[17]), .A2(x[1]), .ZN(n_0_237));
   INV_X1 i_0_318 (.A(n_0_239), .ZN(n_0_238));
   NAND2_X1 i_0_319 (.A1(p[21]), .A2(x[5]), .ZN(n_0_239));
   NOR2_X1 i_0_320 (.A1(p[21]), .A2(x[5]), .ZN(n_0_240));
   INV_X1 i_0_321 (.A(n_0_242), .ZN(n_0_241));
   NAND2_X1 i_0_322 (.A1(p[23]), .A2(x[7]), .ZN(n_0_242));
   NOR2_X1 i_0_323 (.A1(p[23]), .A2(x[7]), .ZN(n_0_243));
   INV_X1 i_0_324 (.A(n_0_245), .ZN(n_0_244));
   NAND2_X1 i_0_325 (.A1(p[25]), .A2(x[9]), .ZN(n_0_245));
   NOR2_X1 i_0_326 (.A1(p[25]), .A2(x[9]), .ZN(n_0_246));
   INV_X1 i_0_327 (.A(n_0_248), .ZN(n_0_247));
   NAND2_X1 i_0_328 (.A1(p[27]), .A2(x[11]), .ZN(n_0_248));
   NOR2_X1 i_0_329 (.A1(p[27]), .A2(x[11]), .ZN(n_0_249));
   INV_X1 i_0_330 (.A(n_0_251), .ZN(n_0_250));
   NAND2_X1 i_0_331 (.A1(p[29]), .A2(x[13]), .ZN(n_0_251));
   NOR2_X1 i_0_332 (.A1(p[29]), .A2(x[13]), .ZN(n_0_252));
   NAND2_X1 i_0_333 (.A1(n_0_257), .A2(i[4]), .ZN(n_120));
   INV_X1 i_0_334 (.A(a[3]), .ZN(n_0_253));
   INV_X1 i_0_335 (.A(a[4]), .ZN(n_0_254));
   INV_X1 i_0_336 (.A(a[8]), .ZN(n_0_255));
   INV_X1 i_0_337 (.A(a[13]), .ZN(n_0_256));
   INV_X1 i_0_338 (.A(reset), .ZN(n_0_257));
   INV_X1 i_0_339 (.A(p[20]), .ZN(n_0_258));
   INV_X1 i_0_340 (.A(i[4]), .ZN(n_0_259));
   INV_X1 i_0_341 (.A(b[8]), .ZN(n_0_260));
   INV_X1 i_0_342 (.A(b[15]), .ZN(n_0_261));
   INV_X1 i_0_343 (.A(n_0_194), .ZN(n_0_262));
   INV_X1 i_0_344 (.A(n_0_193), .ZN(n_0_263));
   INV_X1 i_0_345 (.A(n_0_24), .ZN(n_0_264));
endmodule

module datapath__0_26(result, p_0);
   input [31:0]result;
   output [31:0]p_0;

   HA_X1 i_0 (.A(result[8]), .B(result[7]), .CO(n_0), .S(p_0[8]));
   HA_X1 i_1 (.A(result[9]), .B(n_0), .CO(n_1), .S(p_0[9]));
   HA_X1 i_2 (.A(result[10]), .B(n_1), .CO(n_2), .S(p_0[10]));
   HA_X1 i_3 (.A(result[11]), .B(n_2), .CO(n_3), .S(p_0[11]));
   HA_X1 i_4 (.A(result[12]), .B(n_3), .CO(n_4), .S(p_0[12]));
   HA_X1 i_5 (.A(result[13]), .B(n_4), .CO(n_5), .S(p_0[13]));
   HA_X1 i_6 (.A(result[14]), .B(n_5), .CO(n_6), .S(p_0[14]));
   HA_X1 i_7 (.A(result[15]), .B(n_6), .CO(n_7), .S(p_0[15]));
   HA_X1 i_8 (.A(result[16]), .B(n_7), .CO(n_8), .S(p_0[16]));
   HA_X1 i_9 (.A(result[17]), .B(n_8), .CO(n_9), .S(p_0[17]));
   HA_X1 i_10 (.A(result[18]), .B(n_9), .CO(n_10), .S(p_0[18]));
   HA_X1 i_11 (.A(result[19]), .B(n_10), .CO(n_11), .S(p_0[19]));
   HA_X1 i_12 (.A(result[20]), .B(n_11), .CO(n_12), .S(p_0[20]));
   HA_X1 i_13 (.A(result[21]), .B(n_12), .CO(n_13), .S(p_0[21]));
   HA_X1 i_14 (.A(result[22]), .B(n_13), .CO(n_14), .S(p_0[22]));
   HA_X1 i_15 (.A(result[23]), .B(n_14), .CO(n_15), .S(p_0[23]));
endmodule

module multiplier(multiplicand, multiplier, o_result, overflow_flag, clk, reset);
   input [15:0]multiplicand;
   input [15:0]multiplier;
   output [15:0]o_result;
   output overflow_flag;
   input clk;
   input reset;

   wire [31:0]result;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_1_2;
   wire n_0_1_3;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_1_10;

   shiftadd s (.p(result), .a(multiplicand), .b(multiplier), .clk(clk), .reset(
      reset));
   datapath__0_26 i_0_0 (.result({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, 
      result[23], result[22], result[21], result[20], result[19], result[18], 
      result[17], result[16], result[15], result[14], result[13], result[12], 
      result[11], result[10], result[9], result[8], result[7], uc_8, uc_9, uc_10, 
      uc_11, uc_12, uc_13, uc_14}), .p_0({uc_15, uc_16, uc_17, uc_18, uc_19, 
      uc_20, uc_21, uc_22, o_result[15], o_result[14], o_result[13], 
      o_result[12], o_result[11], o_result[10], o_result[9], o_result[8], 
      o_result[7], o_result[6], o_result[5], o_result[4], o_result[3], 
      o_result[2], o_result[1], o_result[0], uc_23, uc_24, uc_25, uc_26, uc_27, 
      uc_28, uc_29, uc_30}));
   NOR4_X1 i_0_1_0 (.A1(result[0]), .A2(result[1]), .A3(result[2]), .A4(
      result[3]), .ZN(n_0_1_0));
   NOR4_X1 i_0_1_1 (.A1(result[4]), .A2(result[5]), .A3(result[6]), .A4(
      result[7]), .ZN(n_0_1_1));
   NAND2_X1 i_0_1_2 (.A1(n_0_1_0), .A2(n_0_1_1), .ZN(n_0_1_2));
   NAND4_X1 i_0_1_3 (.A1(n_0_1_2), .A2(result[8]), .A3(result[9]), .A4(
      result[10]), .ZN(n_0_1_3));
   NAND4_X1 i_0_1_4 (.A1(result[11]), .A2(result[12]), .A3(result[13]), .A4(
      result[14]), .ZN(n_0_1_4));
   NAND4_X1 i_0_1_5 (.A1(result[15]), .A2(result[16]), .A3(result[17]), .A4(
      result[18]), .ZN(n_0_1_5));
   NAND4_X1 i_0_1_6 (.A1(result[19]), .A2(result[20]), .A3(result[21]), .A4(
      result[22]), .ZN(n_0_1_6));
   NOR4_X1 i_0_1_7 (.A1(n_0_1_3), .A2(n_0_1_4), .A3(n_0_1_5), .A4(n_0_1_6), 
      .ZN(n_0_1_7));
   NOR2_X1 i_0_1_8 (.A1(n_0_1_7), .A2(result[23]), .ZN(n_0_1_8));
   NOR4_X1 i_0_1_9 (.A1(result[24]), .A2(result[25]), .A3(result[26]), .A4(
      result[27]), .ZN(n_0_1_9));
   NOR4_X1 i_0_1_10 (.A1(result[28]), .A2(result[29]), .A3(result[30]), .A4(
      result[31]), .ZN(n_0_1_10));
   NAND3_X1 i_0_1_11 (.A1(n_0_1_8), .A2(n_0_1_9), .A3(n_0_1_10), .ZN(
      overflow_flag));
endmodule
